module hexdecoder(      input [3:0] in,
                        output logic [6:0] out);

// Your code here!


endmodule
