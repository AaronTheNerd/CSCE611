module testtop;

endmodule
